module counter #(
    parameter WIDTH = 8
)(
    //interface signals
    input  logic                 clk,   //clock
    input  logic                 rst, //reset
    input  logic                 en,    // counter enable
    output logic [WIDTH-1:0]     count  // counter output
);

always_ff @(posedge clk or posedge rst)
    if (rst) count <= {WIDTH{1'b0}}; // concatenation to form WIDTH bits of zeros
    else     count <= count + {{WIDTH -1{1'b0}}, en}; // concatenation to form WIDTH-1 bits of 0 and 1 bit of en

endmodule
